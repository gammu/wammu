Wammu
=====

GUI för `Gammu-biblioteket <https://wammu.eu/gammu/>`_.

.. bild:: https://hosted.weblate.org/widgets/gammu/-/svg-badge.svg
    :alt: Översättningsstatus :target:
    https://hosted.weblate.org/engage/gammu/?utm_source=widget

.. bild:: https://landscape.io/github/gammu/wammu/master/landscape.svg?style=flat
    :target: https://landscape.io/github/gammu/wammu/master :alt: Kodhälsa

.. bild:: https://img.shields.io/gratipay/Gammu.svg
    :alt: Gratipay :target: https://gratipay.com/Gammu/

.. bild:: https://www.bountysource.com/badge/team?team_id=23177&style=bounties_received
    :alt: Bountysource :target:
    https://www.bountysource.com/teams/gammu/issues?utm_source=Gammu&utm_medium=shield&utm_campaign=bounties_received

.. bild:: https://travis-ci.org/gammu/wammu.svg?branch=master
    :target: https://travis-ci.org/gammu/wammu

Hemsida
=======

<https://wammu.eu/>

Licens
======

GNU GPL version 3 eller senare.

Första starten
==============

Vid den första starten kommer du att tillfrågas om att ställa in
telefonparametrar. Om du inte använt Gammu/Wammu tidigare kommer
telefonsökning att föreslås, vilket bör lösa problemet för dig.

Användning
==========

Först måste du ansluta till telefonen, sedan kan du utföra åtgärder på
den. För att skapa poster och importera behöver du inte läsa saker från
telefonen, för andra måste du (förvånande? :-)).

Alla åtgärder med aktuell lista är tillgänglig från snabbmenyn för varje
objekt, du kan också använda nycklar: Retur för att redigera och Delete för
att ta bort.

Säkerhetskopiera i huvudmenyn skapar säkerhetskopior på de poster du redan
har hämtat från telefonen.

Felrapportering
===============

Rapportera hittade fel till <https://github.com/gammu/wammu/issues/>.

Översätta
=========

Du kan hjälpa till med att översätta Wammu till ditt språk på
översättningsservern - <https://hosted.weblate.org/projects/gammu/wammu/>.

Versionshantering
=================

Utvecklingen använder Git, huvudgrenen för utveckling är
<git://github.com/gammu/wammu.git>, du kan blädda igenom den via
<https://github.com/gammu/wammu>.
